* Resistors
* Positive to negative -> Smaller knot to bigger numbered knot

V0 OUT 0 0

* Independent Power Sources
VS  VIN 	VOUT 	sin 0 100 50

DA1 VIN  	IN	my-diode
DA2 OUT  	VOUT	my-diode
DA3 VOUT 	IN	my-diode
DA4 OUT  	VIN	my-diode

C1 IN 		OUT 	1u
R2 IN 		OUT 	10k


.MODEL my-diode D

.endc
