* Resistors
* Positive to negative -> Smaller knot to bigger numbered knot

V0 OUT 0 0

* Independent Power Sources
VS  VIN 	VOUT 	sin 0 130.8317 50

DA1 VIN  	IN	my-diode
DA2 OUT  	VOUT	my-diode
DA3 VOUT 	IN	my-diode
DA4 OUT  	VIN	my-diode

* Envelope
*C1 IN 		OUT 	125u
R1 IN 		OUT 	62.5k

.MODEL my-diode D

