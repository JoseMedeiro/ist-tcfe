* Resistors
* Positive to negative -> Smaller knot to bigger numbered knot

R1 1 3 10k

* Independent Power Sources

VS 1 0 sin 10 0.2 50


* Linear dependent Sources

* Diode

DR1 3 0 my-diode

* Test
* V3 4 0 0

.MODEL my-diode D
