* Resistors
* Positive to negative -> Smaller knot to bigger numbered knot

V0 OUT 0 0


* Independent Power Sources
VS  VIN 	VOUT sin 0 130.8317 50


DA1 VIN  	IN	my-diode
DA2 OUT  	VOUT	my-diode
DA3 VOUT 	IN	my-diode
DA4 OUT  	VIN	my-diode

* Envelope
C1 IN 		OUT 	150u
R1 IN 		OUT 	75k


* Diode
R2 	IN 	3 	75k

DR1 3 4 my-diode
DR2 4 5 my-diode
DR3 5 6 my-diode
DR4 6 7 my-diode
DR5 7 8 my-diode
DR6 8 9 my-diode

DR7  9  10 my-diode
DR8  10 11 my-diode
DR9  11 12 my-diode
DR10 12 13 my-diode
DR11 13 14 my-diode
DR12 14 15 my-diode

DR13 15 16 my-diode
DR14 16 17 my-diode
DR15 17 18 my-diode
DR16 18 19 my-diode

DR17 19 20 my-diode
DR18 20 OUT my-diode


* Test
* V3 4 0 0

.MODEL my-diode D

